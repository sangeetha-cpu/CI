�c�                                                                                        �       �����t��pt���y|  1��؎м  ��d|<�t��R��t��}��|�A��U�ZRr=��U�u7��t21��D@�D��D� f�\|f�\f�`|f�\�D p�B�r� p�v��sZ���� ��}� f�ƈd�@f�D�������@�D����f�f�`|f	�uNf�\|f1�f�4��1�f�t;D}7����0������Z�ƻ p��1۸�r��`� ��1�� �����a�&Z|��}���}�4 ��}�. ���GRUB  Geom Hard Disk Read  Error
 � ���< u��         ����   ���                                                U�